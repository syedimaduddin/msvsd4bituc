MACRO FUNCTION
  ORIGIN 0 0 ;
  FOREIGN FUNCTION 0 0 ;
  SIZE 29.24 BY 7.56 ;
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 10.58 4.48 11.78 4.76 ;
      LAYER M2 ;
        RECT 21.76 4.48 22.96 4.76 ;
      LAYER M2 ;
        RECT 11.61 4.48 14.19 4.76 ;
      LAYER M1 ;
        RECT 14.065 4.2 14.315 4.62 ;
      LAYER M2 ;
        RECT 14.19 4.06 21.07 4.34 ;
      LAYER M1 ;
        RECT 20.945 4.2 21.195 4.62 ;
      LAYER M2 ;
        RECT 21.07 4.48 21.93 4.76 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 11.44 4.9 12.64 5.18 ;
      LAYER M2 ;
        RECT 1.12 4.48 2.32 4.76 ;
      LAYER M2 ;
        RECT 9.46 4.9 11.61 5.18 ;
      LAYER M1 ;
        RECT 9.335 4.2 9.585 5.04 ;
      LAYER M2 ;
        RECT 2.58 4.06 9.46 4.34 ;
      LAYER M1 ;
        RECT 2.455 4.2 2.705 4.62 ;
      LAYER M2 ;
        RECT 2.15 4.48 2.58 4.76 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 6.58 4.9 6.86 ;
      LAYER M2 ;
        RECT 8 6.58 9.2 6.86 ;
      LAYER M2 ;
        RECT 14.88 6.58 16.08 6.86 ;
      LAYER M2 ;
        RECT 19.18 6.58 20.38 6.86 ;
      LAYER M3 ;
        RECT 12.76 1.1 13.04 6.88 ;
      LAYER M2 ;
        RECT 4.73 6.58 5.59 6.86 ;
      LAYER M1 ;
        RECT 5.465 6.3 5.715 6.72 ;
      LAYER M2 ;
        RECT 5.59 6.16 8.17 6.44 ;
      LAYER M1 ;
        RECT 8.045 6.3 8.295 6.72 ;
      LAYER M2 ;
        RECT 8.01 6.58 8.33 6.86 ;
      LAYER M2 ;
        RECT 8.17 6.16 13.76 6.44 ;
      LAYER M1 ;
        RECT 13.635 6.3 13.885 6.72 ;
      LAYER M2 ;
        RECT 13.76 6.58 15.05 6.86 ;
      LAYER M2 ;
        RECT 15.75 6.58 16.07 6.86 ;
      LAYER M1 ;
        RECT 15.785 6.3 16.035 6.72 ;
      LAYER M2 ;
        RECT 15.91 6.16 18.49 6.44 ;
      LAYER M1 ;
        RECT 18.365 6.3 18.615 6.72 ;
      LAYER M2 ;
        RECT 18.49 6.58 19.35 6.86 ;
      LAYER M2 ;
        RECT 12.74 6.16 13.06 6.44 ;
      LAYER M3 ;
        RECT 12.76 6.115 13.04 6.485 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.72 0.68 1 6.88 ;
      LAYER M2 ;
        RECT 6.28 6.58 7.48 6.86 ;
      LAYER M2 ;
        RECT 16.6 6.58 17.8 6.86 ;
      LAYER M3 ;
        RECT 25.66 0.68 25.94 6.88 ;
      LAYER M3 ;
        RECT 27.38 0.68 27.66 6.88 ;
      LAYER M3 ;
        RECT 0.72 6.115 1 6.485 ;
      LAYER M4 ;
        RECT 0.86 5.9 6.45 6.7 ;
      LAYER M3 ;
        RECT 6.31 6.3 6.59 6.72 ;
      LAYER M2 ;
        RECT 6.29 6.58 6.61 6.86 ;
      LAYER M4 ;
        RECT 6.45 5.9 16.77 6.7 ;
      LAYER M3 ;
        RECT 16.63 6.3 16.91 6.72 ;
      LAYER M2 ;
        RECT 16.61 6.58 16.93 6.86 ;
      LAYER M4 ;
        RECT 16.77 5.9 25.8 6.7 ;
      LAYER M3 ;
        RECT 25.66 6.115 25.94 6.485 ;
      LAYER M4 ;
        RECT 25.8 5.9 27.52 6.7 ;
      LAYER M3 ;
        RECT 27.38 6.115 27.66 6.485 ;
    END
  END GND
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 19.18 4.48 20.38 4.76 ;
      LAYER M2 ;
        RECT 24.34 4.48 25.54 4.76 ;
      LAYER M2 ;
        RECT 20.05 4.48 20.37 4.76 ;
      LAYER M3 ;
        RECT 20.07 4.62 20.35 5.04 ;
      LAYER M2 ;
        RECT 20.21 4.9 23.65 5.18 ;
      LAYER M1 ;
        RECT 23.525 4.62 23.775 5.04 ;
      LAYER M2 ;
        RECT 23.65 4.48 24.51 4.76 ;
    END
  END D
  PIN F
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 27.78 4.48 28.98 4.76 ;
      LAYER M2 ;
        RECT 14.88 4.48 16.08 4.76 ;
      LAYER M2 ;
        RECT 26.23 4.48 27.95 4.76 ;
      LAYER M1 ;
        RECT 26.105 4.62 26.355 5.04 ;
      LAYER M2 ;
        RECT 24.51 4.9 26.23 5.18 ;
      LAYER M3 ;
        RECT 24.37 4.919 24.65 5.161 ;
      LAYER M4 ;
        RECT 15.91 4.64 24.51 5.44 ;
      LAYER M3 ;
        RECT 15.77 4.62 16.05 5.04 ;
      LAYER M2 ;
        RECT 15.75 4.48 16.07 4.76 ;
    END
  END F
  PIN FN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 6.28 0.28 7.48 0.56 ;
      LAYER M2 ;
        RECT 8 0.28 9.2 0.56 ;
      LAYER M2 ;
        RECT 14.88 0.28 16.08 0.56 ;
      LAYER M2 ;
        RECT 16.6 0.28 17.8 0.56 ;
      LAYER M2 ;
        RECT 21.76 0.28 22.96 0.56 ;
      LAYER M2 ;
        RECT 7.15 0.28 7.47 0.56 ;
      LAYER M3 ;
        RECT 7.17 0 7.45 0.42 ;
      LAYER M4 ;
        RECT 7.31 -0.4 8.17 0.4 ;
      LAYER M3 ;
        RECT 8.03 0 8.31 0.42 ;
      LAYER M2 ;
        RECT 8.01 0.28 8.33 0.56 ;
      LAYER M4 ;
        RECT 8.17 -0.4 14.19 0.4 ;
      LAYER M3 ;
        RECT 14.05 0 14.33 0.42 ;
      LAYER M2 ;
        RECT 14.19 0.28 15.05 0.56 ;
      LAYER M2 ;
        RECT 15.91 0.28 16.77 0.56 ;
      LAYER M2 ;
        RECT 17.47 0.28 17.79 0.56 ;
      LAYER M3 ;
        RECT 17.49 0.42 17.77 1.68 ;
      LAYER M2 ;
        RECT 17.63 1.54 21.07 1.82 ;
      LAYER M1 ;
        RECT 20.945 0.42 21.195 1.68 ;
      LAYER M2 ;
        RECT 21.07 0.28 21.93 0.56 ;
    END
  END FN
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 4.48 4.9 4.76 ;
      LAYER M2 ;
        RECT 6.28 4.48 7.48 4.76 ;
      LAYER M2 ;
        RECT 4.73 4.48 6.45 4.76 ;
    END
  END C
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 16.6 4.48 17.8 4.76 ;
      LAYER M2 ;
        RECT 8 4.48 9.2 4.76 ;
      LAYER M2 ;
        RECT 16.61 4.48 16.93 4.76 ;
      LAYER M1 ;
        RECT 16.645 4.62 16.895 5.04 ;
      LAYER M2 ;
        RECT 13.33 4.9 16.77 5.18 ;
      LAYER M3 ;
        RECT 13.19 4.919 13.47 5.161 ;
      LAYER M4 ;
        RECT 9.89 4.64 13.33 5.44 ;
      LAYER M3 ;
        RECT 9.75 4.62 10.03 5.04 ;
      LAYER M2 ;
        RECT 9.03 4.48 9.89 4.76 ;
    END
  END E
  OBS 
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 10.58 0.28 11.78 0.56 ;
  LAYER M2 ;
        RECT 4.3 0.7 5.16 0.98 ;
  LAYER M1 ;
        RECT 5.035 0 5.285 0.84 ;
  LAYER M2 ;
        RECT 5.16 -0.14 9.89 0.14 ;
  LAYER M1 ;
        RECT 9.765 0 10.015 0.42 ;
  LAYER M2 ;
        RECT 9.89 0.28 10.75 0.56 ;
  LAYER M1 ;
        RECT 5.035 -0.085 5.285 0.085 ;
  LAYER M2 ;
        RECT 4.99 -0.14 5.33 0.14 ;
  LAYER M1 ;
        RECT 5.035 0.755 5.285 0.925 ;
  LAYER M2 ;
        RECT 4.99 0.7 5.33 0.98 ;
  LAYER M1 ;
        RECT 9.765 -0.085 10.015 0.085 ;
  LAYER M2 ;
        RECT 9.72 -0.14 10.06 0.14 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 0.505 ;
  LAYER M2 ;
        RECT 9.72 0.28 10.06 0.56 ;
  LAYER M1 ;
        RECT 5.035 -0.085 5.285 0.085 ;
  LAYER M2 ;
        RECT 4.99 -0.14 5.33 0.14 ;
  LAYER M1 ;
        RECT 5.035 0.755 5.285 0.925 ;
  LAYER M2 ;
        RECT 4.99 0.7 5.33 0.98 ;
  LAYER M1 ;
        RECT 9.765 -0.085 10.015 0.085 ;
  LAYER M2 ;
        RECT 9.72 -0.14 10.06 0.14 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 0.505 ;
  LAYER M2 ;
        RECT 9.72 0.28 10.06 0.56 ;
  LAYER M2 ;
        RECT 19.61 0.7 20.81 0.98 ;
  LAYER M2 ;
        RECT 11.44 0.7 12.64 0.98 ;
  LAYER M2 ;
        RECT 18.92 0.7 19.78 0.98 ;
  LAYER M1 ;
        RECT 18.795 0.84 19.045 1.26 ;
  LAYER M2 ;
        RECT 18.49 1.12 18.92 1.4 ;
  LAYER M1 ;
        RECT 18.365 0 18.615 1.26 ;
  LAYER M2 ;
        RECT 13.76 -0.14 18.49 0.14 ;
  LAYER M1 ;
        RECT 13.635 0 13.885 0.84 ;
  LAYER M2 ;
        RECT 12.47 0.7 13.76 0.98 ;
  LAYER M1 ;
        RECT 13.635 -0.085 13.885 0.085 ;
  LAYER M2 ;
        RECT 13.59 -0.14 13.93 0.14 ;
  LAYER M1 ;
        RECT 13.635 0.755 13.885 0.925 ;
  LAYER M2 ;
        RECT 13.59 0.7 13.93 0.98 ;
  LAYER M1 ;
        RECT 18.365 -0.085 18.615 0.085 ;
  LAYER M2 ;
        RECT 18.32 -0.14 18.66 0.14 ;
  LAYER M1 ;
        RECT 18.365 1.175 18.615 1.345 ;
  LAYER M2 ;
        RECT 18.32 1.12 18.66 1.4 ;
  LAYER M1 ;
        RECT 18.795 0.755 19.045 0.925 ;
  LAYER M2 ;
        RECT 18.75 0.7 19.09 0.98 ;
  LAYER M1 ;
        RECT 18.795 1.175 19.045 1.345 ;
  LAYER M2 ;
        RECT 18.75 1.12 19.09 1.4 ;
  LAYER M1 ;
        RECT 13.635 -0.085 13.885 0.085 ;
  LAYER M2 ;
        RECT 13.59 -0.14 13.93 0.14 ;
  LAYER M1 ;
        RECT 13.635 0.755 13.885 0.925 ;
  LAYER M2 ;
        RECT 13.59 0.7 13.93 0.98 ;
  LAYER M1 ;
        RECT 18.365 -0.085 18.615 0.085 ;
  LAYER M2 ;
        RECT 18.32 -0.14 18.66 0.14 ;
  LAYER M1 ;
        RECT 18.365 1.175 18.615 1.345 ;
  LAYER M2 ;
        RECT 18.32 1.12 18.66 1.4 ;
  LAYER M1 ;
        RECT 18.795 0.755 19.045 0.925 ;
  LAYER M2 ;
        RECT 18.75 0.7 19.09 0.98 ;
  LAYER M1 ;
        RECT 18.795 1.175 19.045 1.345 ;
  LAYER M2 ;
        RECT 18.75 1.12 19.09 1.4 ;
  LAYER M2 ;
        RECT 1.12 0.28 2.32 0.56 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M2 ;
        RECT 24.34 0.28 25.54 0.56 ;
  LAYER M3 ;
        RECT 23.08 0.68 23.36 6.88 ;
  LAYER M2 ;
        RECT 2.15 0.28 3.01 0.56 ;
  LAYER M1 ;
        RECT 2.885 0.42 3.135 1.26 ;
  LAYER M2 ;
        RECT 3.01 1.12 6.02 1.4 ;
  LAYER M3 ;
        RECT 5.88 0.84 6.16 1.26 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M2 ;
        RECT 6.88 0.7 7.74 0.98 ;
  LAYER M3 ;
        RECT 7.6 0.84 7.88 1.26 ;
  LAYER M4 ;
        RECT 7.74 0.86 23.65 1.66 ;
  LAYER M3 ;
        RECT 23.51 0.42 23.79 1.26 ;
  LAYER M2 ;
        RECT 23.65 0.28 24.51 0.56 ;
  LAYER M4 ;
        RECT 23.055 0.86 23.385 1.66 ;
  LAYER M3 ;
        RECT 23.08 1.075 23.36 1.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 0.505 ;
  LAYER M2 ;
        RECT 2.84 0.28 3.18 0.56 ;
  LAYER M1 ;
        RECT 2.885 1.175 3.135 1.345 ;
  LAYER M2 ;
        RECT 2.84 1.12 3.18 1.4 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 0.505 ;
  LAYER M2 ;
        RECT 2.84 0.28 3.18 0.56 ;
  LAYER M1 ;
        RECT 2.885 1.175 3.135 1.345 ;
  LAYER M2 ;
        RECT 2.84 1.12 3.18 1.4 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 0.505 ;
  LAYER M2 ;
        RECT 2.84 0.28 3.18 0.56 ;
  LAYER M1 ;
        RECT 2.885 1.175 3.135 1.345 ;
  LAYER M2 ;
        RECT 2.84 1.12 3.18 1.4 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M2 ;
        RECT 7.58 0.7 7.9 0.98 ;
  LAYER M3 ;
        RECT 7.6 0.68 7.88 1 ;
  LAYER M2 ;
        RECT 23.49 0.28 23.81 0.56 ;
  LAYER M3 ;
        RECT 23.51 0.26 23.79 0.58 ;
  LAYER M3 ;
        RECT 7.6 1.075 7.88 1.445 ;
  LAYER M4 ;
        RECT 7.575 0.86 7.905 1.66 ;
  LAYER M3 ;
        RECT 23.51 1.075 23.79 1.445 ;
  LAYER M4 ;
        RECT 23.485 0.86 23.815 1.66 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 0.505 ;
  LAYER M2 ;
        RECT 2.84 0.28 3.18 0.56 ;
  LAYER M1 ;
        RECT 2.885 1.175 3.135 1.345 ;
  LAYER M2 ;
        RECT 2.84 1.12 3.18 1.4 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M2 ;
        RECT 7.58 0.7 7.9 0.98 ;
  LAYER M3 ;
        RECT 7.6 0.68 7.88 1 ;
  LAYER M2 ;
        RECT 23.49 0.28 23.81 0.56 ;
  LAYER M3 ;
        RECT 23.51 0.26 23.79 0.58 ;
  LAYER M3 ;
        RECT 7.6 1.075 7.88 1.445 ;
  LAYER M4 ;
        RECT 7.575 0.86 7.905 1.66 ;
  LAYER M3 ;
        RECT 23.51 1.075 23.79 1.445 ;
  LAYER M4 ;
        RECT 23.485 0.86 23.815 1.66 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 0.505 ;
  LAYER M2 ;
        RECT 2.84 0.28 3.18 0.56 ;
  LAYER M1 ;
        RECT 2.885 1.175 3.135 1.345 ;
  LAYER M2 ;
        RECT 2.84 1.12 3.18 1.4 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M2 ;
        RECT 7.58 0.7 7.9 0.98 ;
  LAYER M3 ;
        RECT 7.6 0.68 7.88 1 ;
  LAYER M2 ;
        RECT 23.49 0.28 23.81 0.56 ;
  LAYER M3 ;
        RECT 23.51 0.26 23.79 0.58 ;
  LAYER M3 ;
        RECT 7.6 1.075 7.88 1.445 ;
  LAYER M4 ;
        RECT 7.575 0.86 7.905 1.66 ;
  LAYER M3 ;
        RECT 23.08 1.075 23.36 1.445 ;
  LAYER M4 ;
        RECT 23.055 0.86 23.385 1.66 ;
  LAYER M3 ;
        RECT 23.51 1.075 23.79 1.445 ;
  LAYER M4 ;
        RECT 23.485 0.86 23.815 1.66 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 0.505 ;
  LAYER M2 ;
        RECT 2.84 0.28 3.18 0.56 ;
  LAYER M1 ;
        RECT 2.885 1.175 3.135 1.345 ;
  LAYER M2 ;
        RECT 2.84 1.12 3.18 1.4 ;
  LAYER M2 ;
        RECT 5.86 0.7 6.18 0.98 ;
  LAYER M3 ;
        RECT 5.88 0.68 6.16 1 ;
  LAYER M2 ;
        RECT 5.86 1.12 6.18 1.4 ;
  LAYER M3 ;
        RECT 5.88 1.1 6.16 1.42 ;
  LAYER M2 ;
        RECT 7.58 0.7 7.9 0.98 ;
  LAYER M3 ;
        RECT 7.6 0.68 7.88 1 ;
  LAYER M2 ;
        RECT 23.49 0.28 23.81 0.56 ;
  LAYER M3 ;
        RECT 23.51 0.26 23.79 0.58 ;
  LAYER M3 ;
        RECT 7.6 1.075 7.88 1.445 ;
  LAYER M4 ;
        RECT 7.575 0.86 7.905 1.66 ;
  LAYER M3 ;
        RECT 23.08 1.075 23.36 1.445 ;
  LAYER M4 ;
        RECT 23.055 0.86 23.385 1.66 ;
  LAYER M3 ;
        RECT 23.51 1.075 23.79 1.445 ;
  LAYER M4 ;
        RECT 23.485 0.86 23.815 1.66 ;
  LAYER M2 ;
        RECT 17.03 0.7 18.23 0.98 ;
  LAYER M2 ;
        RECT 27.78 0.28 28.98 0.56 ;
  LAYER M2 ;
        RECT 17.9 0.7 18.22 0.98 ;
  LAYER M3 ;
        RECT 17.92 0 18.2 0.84 ;
  LAYER M4 ;
        RECT 18.06 -0.4 26.23 0.4 ;
  LAYER M3 ;
        RECT 26.09 0 26.37 0.42 ;
  LAYER M2 ;
        RECT 26.23 0.28 27.95 0.56 ;
  LAYER M2 ;
        RECT 17.9 0.7 18.22 0.98 ;
  LAYER M3 ;
        RECT 17.92 0.68 18.2 1 ;
  LAYER M2 ;
        RECT 26.07 0.28 26.39 0.56 ;
  LAYER M3 ;
        RECT 26.09 0.26 26.37 0.58 ;
  LAYER M3 ;
        RECT 17.92 -0.185 18.2 0.185 ;
  LAYER M4 ;
        RECT 17.895 -0.4 18.225 0.4 ;
  LAYER M3 ;
        RECT 26.09 -0.185 26.37 0.185 ;
  LAYER M4 ;
        RECT 26.065 -0.4 26.395 0.4 ;
  LAYER M2 ;
        RECT 17.9 0.7 18.22 0.98 ;
  LAYER M3 ;
        RECT 17.92 0.68 18.2 1 ;
  LAYER M2 ;
        RECT 26.07 0.28 26.39 0.56 ;
  LAYER M3 ;
        RECT 26.09 0.26 26.37 0.58 ;
  LAYER M3 ;
        RECT 17.92 -0.185 18.2 0.185 ;
  LAYER M4 ;
        RECT 17.895 -0.4 18.225 0.4 ;
  LAYER M3 ;
        RECT 26.09 -0.185 26.37 0.185 ;
  LAYER M4 ;
        RECT 26.065 -0.4 26.395 0.4 ;
  LAYER M2 ;
        RECT 3.7 0.28 4.9 0.56 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M2 ;
        RECT 14.45 0.7 15.65 0.98 ;
  LAYER M2 ;
        RECT 19.18 0.28 20.38 0.56 ;
  LAYER M2 ;
        RECT 4.73 0.28 5.59 0.56 ;
  LAYER M3 ;
        RECT 5.45 0.42 5.73 1.26 ;
  LAYER M4 ;
        RECT 5.59 0.86 6.88 1.66 ;
  LAYER M3 ;
        RECT 6.74 1.26 7.02 1.68 ;
  LAYER M2 ;
        RECT 6.88 1.54 8.6 1.82 ;
  LAYER M3 ;
        RECT 8.46 0.84 8.74 1.68 ;
  LAYER M2 ;
        RECT 8.44 0.7 8.76 0.98 ;
  LAYER M2 ;
        RECT 8.6 1.54 14.62 1.82 ;
  LAYER M3 ;
        RECT 14.48 0.84 14.76 1.68 ;
  LAYER M2 ;
        RECT 14.46 0.7 14.78 0.98 ;
  LAYER M3 ;
        RECT 14.48 1.68 14.76 2.1 ;
  LAYER M2 ;
        RECT 14.62 1.96 18.49 2.24 ;
  LAYER M3 ;
        RECT 18.35 0.42 18.63 2.1 ;
  LAYER M2 ;
        RECT 18.49 0.28 19.35 0.56 ;
  LAYER M2 ;
        RECT 5.43 0.28 5.75 0.56 ;
  LAYER M3 ;
        RECT 5.45 0.26 5.73 0.58 ;
  LAYER M2 ;
        RECT 6.72 1.54 7.04 1.82 ;
  LAYER M3 ;
        RECT 6.74 1.52 7.02 1.84 ;
  LAYER M2 ;
        RECT 8.44 0.7 8.76 0.98 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 1 ;
  LAYER M2 ;
        RECT 8.44 1.54 8.76 1.82 ;
  LAYER M3 ;
        RECT 8.46 1.52 8.74 1.84 ;
  LAYER M3 ;
        RECT 5.45 1.075 5.73 1.445 ;
  LAYER M4 ;
        RECT 5.425 0.86 5.755 1.66 ;
  LAYER M3 ;
        RECT 6.74 1.075 7.02 1.445 ;
  LAYER M4 ;
        RECT 6.715 0.86 7.045 1.66 ;
  LAYER M2 ;
        RECT 5.43 0.28 5.75 0.56 ;
  LAYER M3 ;
        RECT 5.45 0.26 5.73 0.58 ;
  LAYER M2 ;
        RECT 6.72 1.54 7.04 1.82 ;
  LAYER M3 ;
        RECT 6.74 1.52 7.02 1.84 ;
  LAYER M2 ;
        RECT 8.44 0.7 8.76 0.98 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 1 ;
  LAYER M2 ;
        RECT 8.44 1.54 8.76 1.82 ;
  LAYER M3 ;
        RECT 8.46 1.52 8.74 1.84 ;
  LAYER M3 ;
        RECT 5.45 1.075 5.73 1.445 ;
  LAYER M4 ;
        RECT 5.425 0.86 5.755 1.66 ;
  LAYER M3 ;
        RECT 6.74 1.075 7.02 1.445 ;
  LAYER M4 ;
        RECT 6.715 0.86 7.045 1.66 ;
  LAYER M2 ;
        RECT 5.43 0.28 5.75 0.56 ;
  LAYER M3 ;
        RECT 5.45 0.26 5.73 0.58 ;
  LAYER M2 ;
        RECT 6.72 1.54 7.04 1.82 ;
  LAYER M3 ;
        RECT 6.74 1.52 7.02 1.84 ;
  LAYER M2 ;
        RECT 8.44 0.7 8.76 0.98 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 1 ;
  LAYER M2 ;
        RECT 8.44 1.54 8.76 1.82 ;
  LAYER M3 ;
        RECT 8.46 1.52 8.74 1.84 ;
  LAYER M2 ;
        RECT 14.46 0.7 14.78 0.98 ;
  LAYER M3 ;
        RECT 14.48 0.68 14.76 1 ;
  LAYER M2 ;
        RECT 14.46 1.54 14.78 1.82 ;
  LAYER M3 ;
        RECT 14.48 1.52 14.76 1.84 ;
  LAYER M3 ;
        RECT 5.45 1.075 5.73 1.445 ;
  LAYER M4 ;
        RECT 5.425 0.86 5.755 1.66 ;
  LAYER M3 ;
        RECT 6.74 1.075 7.02 1.445 ;
  LAYER M4 ;
        RECT 6.715 0.86 7.045 1.66 ;
  LAYER M2 ;
        RECT 5.43 0.28 5.75 0.56 ;
  LAYER M3 ;
        RECT 5.45 0.26 5.73 0.58 ;
  LAYER M2 ;
        RECT 6.72 1.54 7.04 1.82 ;
  LAYER M3 ;
        RECT 6.74 1.52 7.02 1.84 ;
  LAYER M2 ;
        RECT 8.44 0.7 8.76 0.98 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 1 ;
  LAYER M2 ;
        RECT 8.44 1.54 8.76 1.82 ;
  LAYER M3 ;
        RECT 8.46 1.52 8.74 1.84 ;
  LAYER M2 ;
        RECT 14.46 0.7 14.78 0.98 ;
  LAYER M3 ;
        RECT 14.48 0.68 14.76 1 ;
  LAYER M2 ;
        RECT 14.46 1.54 14.78 1.82 ;
  LAYER M3 ;
        RECT 14.48 1.52 14.76 1.84 ;
  LAYER M3 ;
        RECT 5.45 1.075 5.73 1.445 ;
  LAYER M4 ;
        RECT 5.425 0.86 5.755 1.66 ;
  LAYER M3 ;
        RECT 6.74 1.075 7.02 1.445 ;
  LAYER M4 ;
        RECT 6.715 0.86 7.045 1.66 ;
  LAYER M2 ;
        RECT 5.43 0.28 5.75 0.56 ;
  LAYER M3 ;
        RECT 5.45 0.26 5.73 0.58 ;
  LAYER M2 ;
        RECT 6.72 1.54 7.04 1.82 ;
  LAYER M3 ;
        RECT 6.74 1.52 7.02 1.84 ;
  LAYER M2 ;
        RECT 8.44 0.7 8.76 0.98 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 1 ;
  LAYER M2 ;
        RECT 8.44 1.54 8.76 1.82 ;
  LAYER M3 ;
        RECT 8.46 1.52 8.74 1.84 ;
  LAYER M2 ;
        RECT 14.46 0.7 14.78 0.98 ;
  LAYER M3 ;
        RECT 14.48 0.68 14.76 1 ;
  LAYER M2 ;
        RECT 14.46 1.54 14.78 1.82 ;
  LAYER M3 ;
        RECT 14.48 1.52 14.76 1.84 ;
  LAYER M2 ;
        RECT 14.46 1.96 14.78 2.24 ;
  LAYER M3 ;
        RECT 14.48 1.94 14.76 2.26 ;
  LAYER M2 ;
        RECT 18.33 0.28 18.65 0.56 ;
  LAYER M3 ;
        RECT 18.35 0.26 18.63 0.58 ;
  LAYER M2 ;
        RECT 18.33 1.96 18.65 2.24 ;
  LAYER M3 ;
        RECT 18.35 1.94 18.63 2.26 ;
  LAYER M3 ;
        RECT 5.45 1.075 5.73 1.445 ;
  LAYER M4 ;
        RECT 5.425 0.86 5.755 1.66 ;
  LAYER M3 ;
        RECT 6.74 1.075 7.02 1.445 ;
  LAYER M4 ;
        RECT 6.715 0.86 7.045 1.66 ;
  LAYER M2 ;
        RECT 5.43 0.28 5.75 0.56 ;
  LAYER M3 ;
        RECT 5.45 0.26 5.73 0.58 ;
  LAYER M2 ;
        RECT 6.72 1.54 7.04 1.82 ;
  LAYER M3 ;
        RECT 6.74 1.52 7.02 1.84 ;
  LAYER M2 ;
        RECT 8.44 0.7 8.76 0.98 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 1 ;
  LAYER M2 ;
        RECT 8.44 1.54 8.76 1.82 ;
  LAYER M3 ;
        RECT 8.46 1.52 8.74 1.84 ;
  LAYER M2 ;
        RECT 14.46 0.7 14.78 0.98 ;
  LAYER M3 ;
        RECT 14.48 0.68 14.76 1 ;
  LAYER M2 ;
        RECT 14.46 1.54 14.78 1.82 ;
  LAYER M3 ;
        RECT 14.48 1.52 14.76 1.84 ;
  LAYER M2 ;
        RECT 14.46 1.96 14.78 2.24 ;
  LAYER M3 ;
        RECT 14.48 1.94 14.76 2.26 ;
  LAYER M2 ;
        RECT 18.33 0.28 18.65 0.56 ;
  LAYER M3 ;
        RECT 18.35 0.26 18.63 0.58 ;
  LAYER M2 ;
        RECT 18.33 1.96 18.65 2.24 ;
  LAYER M3 ;
        RECT 18.35 1.94 18.63 2.26 ;
  LAYER M3 ;
        RECT 5.45 1.075 5.73 1.445 ;
  LAYER M4 ;
        RECT 5.425 0.86 5.755 1.66 ;
  LAYER M3 ;
        RECT 6.74 1.075 7.02 1.445 ;
  LAYER M4 ;
        RECT 6.715 0.86 7.045 1.66 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 3.865 ;
  LAYER M1 ;
        RECT 11.485 4.115 11.735 5.125 ;
  LAYER M1 ;
        RECT 11.485 6.215 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.055 0.335 11.305 3.865 ;
  LAYER M1 ;
        RECT 11.915 0.335 12.165 3.865 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 3.865 ;
  LAYER M1 ;
        RECT 12.345 4.115 12.595 5.125 ;
  LAYER M1 ;
        RECT 12.345 6.215 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.775 0.335 13.025 3.865 ;
  LAYER M2 ;
        RECT 11.01 1.12 13.07 1.4 ;
  LAYER M2 ;
        RECT 11.44 6.58 13.07 6.86 ;
  LAYER M2 ;
        RECT 10.58 0.28 11.78 0.56 ;
  LAYER M2 ;
        RECT 11.44 0.7 12.64 0.98 ;
  LAYER M2 ;
        RECT 10.58 4.48 11.78 4.76 ;
  LAYER M2 ;
        RECT 11.44 4.9 12.64 5.18 ;
  LAYER M3 ;
        RECT 12.76 1.1 13.04 6.88 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 3.865 ;
  LAYER M1 ;
        RECT 1.165 4.115 1.415 5.125 ;
  LAYER M1 ;
        RECT 1.165 6.215 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.595 0.335 1.845 3.865 ;
  LAYER M1 ;
        RECT 0.735 0.335 0.985 3.865 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.28 2.32 0.56 ;
  LAYER M2 ;
        RECT 1.12 4.48 2.32 4.76 ;
  LAYER M3 ;
        RECT 0.72 0.68 1 6.88 ;
  LAYER M1 ;
        RECT 25.245 0.335 25.495 3.865 ;
  LAYER M1 ;
        RECT 25.245 4.115 25.495 5.125 ;
  LAYER M1 ;
        RECT 25.245 6.215 25.495 7.225 ;
  LAYER M1 ;
        RECT 24.815 0.335 25.065 3.865 ;
  LAYER M1 ;
        RECT 25.675 0.335 25.925 3.865 ;
  LAYER M2 ;
        RECT 24.77 0.7 25.97 0.98 ;
  LAYER M2 ;
        RECT 24.77 6.58 25.97 6.86 ;
  LAYER M2 ;
        RECT 24.34 0.28 25.54 0.56 ;
  LAYER M2 ;
        RECT 24.34 4.48 25.54 4.76 ;
  LAYER M3 ;
        RECT 25.66 0.68 25.94 6.88 ;
  LAYER M1 ;
        RECT 27.825 0.335 28.075 3.865 ;
  LAYER M1 ;
        RECT 27.825 4.115 28.075 5.125 ;
  LAYER M1 ;
        RECT 27.825 6.215 28.075 7.225 ;
  LAYER M1 ;
        RECT 28.255 0.335 28.505 3.865 ;
  LAYER M1 ;
        RECT 27.395 0.335 27.645 3.865 ;
  LAYER M2 ;
        RECT 27.35 0.7 28.55 0.98 ;
  LAYER M2 ;
        RECT 27.35 6.58 28.55 6.86 ;
  LAYER M2 ;
        RECT 27.78 0.28 28.98 0.56 ;
  LAYER M2 ;
        RECT 27.78 4.48 28.98 4.76 ;
  LAYER M3 ;
        RECT 27.38 0.68 27.66 6.88 ;
  LAYER M1 ;
        RECT 22.665 0.335 22.915 3.865 ;
  LAYER M1 ;
        RECT 22.665 4.115 22.915 5.125 ;
  LAYER M1 ;
        RECT 22.665 6.215 22.915 7.225 ;
  LAYER M1 ;
        RECT 22.235 0.335 22.485 3.865 ;
  LAYER M1 ;
        RECT 23.095 0.335 23.345 3.865 ;
  LAYER M2 ;
        RECT 22.19 0.7 23.39 0.98 ;
  LAYER M2 ;
        RECT 22.19 6.58 23.39 6.86 ;
  LAYER M2 ;
        RECT 21.76 0.28 22.96 0.56 ;
  LAYER M2 ;
        RECT 21.76 4.48 22.96 4.76 ;
  LAYER M3 ;
        RECT 23.08 0.68 23.36 6.88 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 3.865 ;
  LAYER M1 ;
        RECT 6.325 4.115 6.575 5.125 ;
  LAYER M1 ;
        RECT 6.325 6.215 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.755 0.335 7.005 3.865 ;
  LAYER M1 ;
        RECT 5.895 0.335 6.145 3.865 ;
  LAYER M2 ;
        RECT 6.28 6.58 7.48 6.86 ;
  LAYER M2 ;
        RECT 6.28 0.28 7.48 0.56 ;
  LAYER M2 ;
        RECT 6.28 4.48 7.48 4.76 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M1 ;
        RECT 17.505 0.335 17.755 3.865 ;
  LAYER M1 ;
        RECT 17.505 4.115 17.755 5.125 ;
  LAYER M1 ;
        RECT 17.505 6.215 17.755 7.225 ;
  LAYER M1 ;
        RECT 17.075 0.335 17.325 3.865 ;
  LAYER M1 ;
        RECT 17.935 0.335 18.185 3.865 ;
  LAYER M2 ;
        RECT 16.6 6.58 17.8 6.86 ;
  LAYER M2 ;
        RECT 16.6 0.28 17.8 0.56 ;
  LAYER M2 ;
        RECT 16.6 4.48 17.8 4.76 ;
  LAYER M2 ;
        RECT 17.03 0.7 18.23 0.98 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 3.865 ;
  LAYER M1 ;
        RECT 3.745 4.115 3.995 5.125 ;
  LAYER M1 ;
        RECT 3.745 6.215 3.995 7.225 ;
  LAYER M1 ;
        RECT 4.175 0.335 4.425 3.865 ;
  LAYER M1 ;
        RECT 3.315 0.335 3.565 3.865 ;
  LAYER M2 ;
        RECT 3.7 6.58 4.9 6.86 ;
  LAYER M2 ;
        RECT 3.7 0.28 4.9 0.56 ;
  LAYER M2 ;
        RECT 3.7 4.48 4.9 4.76 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M1 ;
        RECT 20.085 0.335 20.335 3.865 ;
  LAYER M1 ;
        RECT 20.085 4.115 20.335 5.125 ;
  LAYER M1 ;
        RECT 20.085 6.215 20.335 7.225 ;
  LAYER M1 ;
        RECT 19.655 0.335 19.905 3.865 ;
  LAYER M1 ;
        RECT 20.515 0.335 20.765 3.865 ;
  LAYER M2 ;
        RECT 19.18 6.58 20.38 6.86 ;
  LAYER M2 ;
        RECT 19.18 0.28 20.38 0.56 ;
  LAYER M2 ;
        RECT 19.18 4.48 20.38 4.76 ;
  LAYER M2 ;
        RECT 19.61 0.7 20.81 0.98 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 3.865 ;
  LAYER M1 ;
        RECT 8.905 4.115 9.155 5.125 ;
  LAYER M1 ;
        RECT 8.905 6.215 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.475 0.335 8.725 3.865 ;
  LAYER M1 ;
        RECT 9.335 0.335 9.585 3.865 ;
  LAYER M2 ;
        RECT 8 6.58 9.2 6.86 ;
  LAYER M2 ;
        RECT 8 0.28 9.2 0.56 ;
  LAYER M2 ;
        RECT 8 4.48 9.2 4.76 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 3.865 ;
  LAYER M1 ;
        RECT 14.925 4.115 15.175 5.125 ;
  LAYER M1 ;
        RECT 14.925 6.215 15.175 7.225 ;
  LAYER M1 ;
        RECT 15.355 0.335 15.605 3.865 ;
  LAYER M1 ;
        RECT 14.495 0.335 14.745 3.865 ;
  LAYER M2 ;
        RECT 14.88 6.58 16.08 6.86 ;
  LAYER M2 ;
        RECT 14.88 0.28 16.08 0.56 ;
  LAYER M2 ;
        RECT 14.88 4.48 16.08 4.76 ;
  LAYER M2 ;
        RECT 14.45 0.7 15.65 0.98 ;
  END 
END FUNCTION

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RING_OSCILLATOR
  CLASS BLOCK ;
  FOREIGN RING_OSCILLATOR ;
  ORIGIN 0.590 0.590 ;
  SIZE 13.020 BY 15.710 ;
  PIN VDD
    ANTENNADIFFAREA 3.910200 ;
    PORT
      LAYER nwell ;
        RECT 0.000 7.560 7.740 15.120 ;
      LAYER li1 ;
        RECT 1.165 13.775 1.415 14.785 ;
        RECT 3.745 13.775 3.995 14.785 ;
        RECT 6.325 13.775 6.575 14.785 ;
        RECT 0.735 7.895 0.985 11.425 ;
        RECT 1.595 7.895 1.845 11.425 ;
        RECT 2.885 -0.085 3.135 9.325 ;
        RECT 3.315 7.895 3.565 11.425 ;
        RECT 4.175 7.895 4.425 11.425 ;
        RECT 5.895 7.895 6.145 11.425 ;
        RECT 6.755 7.895 7.005 11.425 ;
        RECT 7.185 -0.085 7.435 8.905 ;
      LAYER mcon ;
        RECT 1.205 14.195 1.375 14.365 ;
        RECT 3.785 14.195 3.955 14.365 ;
        RECT 6.365 14.195 6.535 14.365 ;
        RECT 0.775 8.315 0.945 8.485 ;
        RECT 1.635 8.315 1.805 8.485 ;
        RECT 2.925 9.155 3.095 9.325 ;
        RECT 3.355 8.315 3.525 8.485 ;
        RECT 4.215 8.315 4.385 8.485 ;
        RECT 5.935 8.315 6.105 8.485 ;
        RECT 6.795 8.315 6.965 8.485 ;
        RECT 7.225 8.735 7.395 8.905 ;
        RECT 2.925 -0.085 3.095 0.085 ;
        RECT 7.225 -0.085 7.395 0.085 ;
      LAYER met1 ;
        RECT 0.690 14.140 1.890 14.420 ;
        RECT 3.270 14.140 4.470 14.420 ;
        RECT 5.850 14.140 7.050 14.420 ;
        RECT 2.840 9.100 3.600 9.380 ;
        RECT 0.700 8.680 1.450 8.960 ;
        RECT 6.720 8.680 7.480 8.960 ;
        RECT 0.690 8.260 1.890 8.540 ;
        RECT 3.270 8.260 4.470 8.540 ;
        RECT 5.850 8.260 7.050 8.540 ;
        RECT 2.840 -0.140 3.180 0.140 ;
        RECT 6.290 -0.140 7.480 0.140 ;
      LAYER via ;
        RECT 0.730 14.150 0.990 14.410 ;
        RECT 3.310 14.150 3.570 14.410 ;
        RECT 6.750 14.150 7.010 14.410 ;
        RECT 3.310 9.110 3.570 9.370 ;
        RECT 0.730 8.690 0.990 8.950 ;
        RECT 1.160 8.690 1.420 8.950 ;
        RECT 6.750 8.690 7.010 8.950 ;
        RECT 0.730 8.270 0.990 8.530 ;
        RECT 3.310 8.270 3.570 8.530 ;
        RECT 6.750 8.270 7.010 8.530 ;
        RECT 2.880 -0.130 3.140 0.130 ;
        RECT 6.320 -0.130 6.580 0.130 ;
      LAYER met2 ;
        RECT 0.720 8.240 1.000 14.440 ;
        RECT 1.150 -0.185 1.430 8.980 ;
        RECT 3.300 8.240 3.580 14.440 ;
        RECT 6.740 8.240 7.020 14.440 ;
        RECT 2.870 -0.185 3.150 0.240 ;
        RECT 6.310 -0.185 6.590 0.240 ;
      LAYER via2 ;
        RECT 1.150 -0.140 1.430 0.140 ;
        RECT 2.870 -0.140 3.150 0.140 ;
        RECT 6.310 -0.140 6.590 0.140 ;
      LAYER met3 ;
        RECT -0.400 -0.400 12.240 0.400 ;
      LAYER via3 ;
        RECT -0.160 -0.160 0.160 0.160 ;
      LAYER met4 ;
        RECT -0.590 -0.590 0.590 9.410 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 3.910200 ;
    PORT
      LAYER pwell ;
        RECT 1.075 0.150 1.505 1.530 ;
        RECT 3.655 0.150 4.085 1.530 ;
        RECT 6.235 0.150 6.665 1.530 ;
      LAYER li1 ;
        RECT 0.735 3.695 0.985 7.225 ;
        RECT 1.595 3.695 1.845 7.225 ;
        RECT 3.315 3.695 3.565 7.225 ;
        RECT 4.175 3.695 4.425 7.225 ;
        RECT 5.895 3.695 6.145 7.225 ;
        RECT 6.755 3.695 7.005 7.225 ;
        RECT 1.165 0.335 1.415 1.345 ;
        RECT 3.745 0.335 3.995 1.345 ;
        RECT 6.325 0.335 6.575 1.345 ;
      LAYER mcon ;
        RECT 0.775 6.635 0.945 6.805 ;
        RECT 1.635 6.635 1.805 6.805 ;
        RECT 3.355 6.635 3.525 6.805 ;
        RECT 4.215 6.635 4.385 6.805 ;
        RECT 5.935 6.635 6.105 6.805 ;
        RECT 6.795 6.635 6.965 6.805 ;
        RECT 1.205 0.755 1.375 0.925 ;
        RECT 3.785 0.755 3.955 0.925 ;
        RECT 6.365 0.755 6.535 0.925 ;
      LAYER met1 ;
        RECT 0.690 6.580 1.890 6.860 ;
        RECT 3.270 6.580 4.470 6.860 ;
        RECT 5.850 6.580 7.050 6.860 ;
        RECT 0.270 6.160 1.020 6.440 ;
        RECT 2.850 6.160 3.600 6.440 ;
        RECT 6.290 6.160 7.040 6.440 ;
        RECT 0.690 0.700 1.890 0.980 ;
        RECT 3.270 0.700 4.470 0.980 ;
        RECT 5.850 0.700 7.050 0.980 ;
      LAYER via ;
        RECT 0.730 6.590 0.990 6.850 ;
        RECT 3.310 6.590 3.570 6.850 ;
        RECT 6.750 6.590 7.010 6.850 ;
        RECT 0.300 6.170 0.560 6.430 ;
        RECT 0.730 6.170 0.990 6.430 ;
        RECT 2.880 6.170 3.140 6.430 ;
        RECT 3.310 6.170 3.570 6.430 ;
        RECT 6.320 6.170 6.580 6.430 ;
        RECT 6.750 6.170 7.010 6.430 ;
        RECT 0.730 0.710 0.990 0.970 ;
        RECT 3.310 0.710 3.570 0.970 ;
        RECT 6.750 0.710 7.010 0.970 ;
      LAYER met2 ;
        RECT 0.290 6.140 0.570 9.005 ;
        RECT 0.720 0.680 1.000 6.880 ;
        RECT 2.870 6.140 3.150 9.005 ;
        RECT 3.300 0.680 3.580 6.880 ;
        RECT 6.310 6.140 6.590 9.005 ;
        RECT 6.740 0.680 7.020 6.880 ;
      LAYER via2 ;
        RECT 0.290 8.680 0.570 8.960 ;
        RECT 2.870 8.680 3.150 8.960 ;
        RECT 6.310 8.680 6.590 8.960 ;
      LAYER met3 ;
        RECT -0.400 8.420 12.240 9.220 ;
      LAYER via3 ;
        RECT 11.680 8.660 12.000 8.980 ;
      LAYER met4 ;
        RECT 11.250 -0.590 12.430 9.410 ;
    END
  END VSS
  PIN INP
    ANTENNAGATEAREA 1.260000 ;
    ANTENNADIFFAREA 1.176000 ;
    PORT
      LAYER li1 ;
        RECT 3.745 11.675 3.995 12.685 ;
        RECT 1.165 7.895 1.415 11.425 ;
        RECT 1.165 3.695 1.415 7.225 ;
        RECT 3.745 2.435 3.995 3.445 ;
      LAYER mcon ;
        RECT 3.785 12.095 3.955 12.265 ;
        RECT 1.205 7.895 1.375 8.065 ;
        RECT 1.205 7.055 1.375 7.225 ;
        RECT 3.785 2.855 3.955 3.025 ;
      LAYER met1 ;
        RECT 3.700 12.040 4.900 12.320 ;
        RECT 1.120 7.840 2.320 8.120 ;
        RECT 1.560 7.420 4.460 7.700 ;
        RECT 1.120 7.000 2.320 7.280 ;
        RECT 3.700 2.800 4.900 3.080 ;
      LAYER via ;
        RECT 4.170 12.050 4.430 12.310 ;
        RECT 1.590 7.850 1.850 8.110 ;
        RECT 1.590 7.430 1.850 7.690 ;
        RECT 4.170 7.430 4.430 7.690 ;
        RECT 1.590 7.010 1.850 7.270 ;
        RECT 4.170 2.810 4.430 3.070 ;
      LAYER met2 ;
        RECT 1.580 6.980 1.860 8.140 ;
        RECT 4.160 2.780 4.440 12.340 ;
    END
  END INP
  OBS
      LAYER pwell ;
        RECT 0.605 3.545 1.975 5.905 ;
        RECT 3.185 3.545 4.555 5.905 ;
        RECT 5.765 3.545 7.135 5.905 ;
      LAYER li1 ;
        RECT 1.165 11.675 1.415 12.685 ;
        RECT 1.165 2.435 1.415 3.445 ;
        RECT 2.025 2.855 2.275 12.265 ;
        RECT 3.745 7.895 3.995 11.425 ;
        RECT 3.745 3.695 3.995 7.225 ;
        RECT 4.605 6.215 4.855 11.845 ;
        RECT 5.465 11.675 5.715 12.265 ;
        RECT 6.325 11.675 6.575 12.685 ;
        RECT 6.325 7.895 6.575 11.425 ;
        RECT 5.465 2.855 5.715 6.385 ;
        RECT 6.325 3.695 6.575 7.225 ;
        RECT 6.325 2.435 6.575 3.445 ;
      LAYER mcon ;
        RECT 1.205 12.095 1.375 12.265 ;
        RECT 2.065 12.095 2.235 12.265 ;
        RECT 5.505 12.095 5.675 12.265 ;
        RECT 4.645 11.675 4.815 11.845 ;
        RECT 5.505 11.675 5.675 11.845 ;
        RECT 6.365 12.095 6.535 12.265 ;
        RECT 2.065 8.735 2.235 8.905 ;
        RECT 1.205 2.855 1.375 3.025 ;
        RECT 3.785 7.895 3.955 8.065 ;
        RECT 4.645 7.895 4.815 8.065 ;
        RECT 6.365 7.895 6.535 8.065 ;
        RECT 3.785 7.055 3.955 7.225 ;
        RECT 4.645 7.055 4.815 7.225 ;
        RECT 6.365 7.055 6.535 7.225 ;
        RECT 4.645 6.215 4.815 6.385 ;
        RECT 5.505 6.215 5.675 6.385 ;
        RECT 2.065 2.855 2.235 3.025 ;
        RECT 5.505 2.855 5.675 3.025 ;
        RECT 6.365 2.855 6.535 3.025 ;
      LAYER met1 ;
        RECT 1.120 12.040 2.320 12.320 ;
        RECT 5.420 12.040 6.620 12.320 ;
        RECT 4.560 11.620 5.760 11.900 ;
        RECT 1.980 8.680 5.750 8.960 ;
        RECT 3.700 7.840 4.900 8.120 ;
        RECT 5.420 7.840 6.620 8.120 ;
        RECT 3.700 7.000 4.900 7.280 ;
        RECT 5.420 7.000 6.620 7.280 ;
        RECT 4.560 6.160 5.760 6.440 ;
        RECT 1.120 2.800 2.320 3.080 ;
        RECT 5.420 2.800 6.620 3.080 ;
      LAYER via ;
        RECT 5.460 8.690 5.720 8.950 ;
        RECT 5.460 7.850 5.720 8.110 ;
        RECT 5.890 7.850 6.150 8.110 ;
        RECT 5.890 7.010 6.150 7.270 ;
      LAYER met2 ;
        RECT 5.450 7.820 5.730 8.980 ;
        RECT 5.880 6.980 6.160 8.140 ;
  END
END RING_OSCILLATOR
END LIBRARY


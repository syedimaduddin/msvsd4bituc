module ADC_1BIT(
	output OUT,
	input INN,
	input INP
);

endmodule

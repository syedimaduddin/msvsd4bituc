VERSION 5.7 ;

  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ADC_1BIT
  CLASS BLOCK ;
  FOREIGN ADC_1BIT ;
  ORIGIN -0.260 0.000 ;
  SIZE 10.920 BY 15.280 ;
  PIN VSS
    ANTENNADIFFAREA 3.385200 ;
    PORT
      LAYER pwell ;
        RECT 3.655 0.150 4.945 1.530 ;
        RECT 7.095 0.150 7.525 1.530 ;
      LAYER li1 ;
        RECT 3.315 3.695 3.565 7.225 ;
        RECT 4.175 3.695 4.425 7.225 ;
        RECT 5.035 3.695 5.285 7.225 ;
        RECT 6.755 3.695 7.005 7.225 ;
        RECT 7.615 3.695 7.865 7.225 ;
        RECT 3.745 0.335 3.995 1.345 ;
        RECT 4.605 0.335 4.855 1.345 ;
        RECT 7.185 0.335 7.435 1.345 ;
      LAYER mcon ;
        RECT 3.355 6.215 3.525 6.385 ;
        RECT 4.215 6.215 4.385 6.385 ;
        RECT 5.075 6.215 5.245 6.385 ;
        RECT 6.795 6.635 6.965 6.805 ;
        RECT 7.655 6.635 7.825 6.805 ;
        RECT 3.785 0.755 3.955 0.925 ;
        RECT 4.645 0.755 4.815 0.925 ;
        RECT 7.225 0.755 7.395 0.925 ;
      LAYER met1 ;
        RECT 6.710 6.580 7.910 6.860 ;
        RECT 3.270 6.160 5.330 6.440 ;
        RECT 3.710 3.640 7.040 3.920 ;
        RECT 3.700 0.700 4.900 0.980 ;
        RECT 6.710 0.700 7.910 0.980 ;
      LAYER via ;
        RECT 6.750 6.590 7.010 6.850 ;
        RECT 3.740 6.170 4.000 6.430 ;
        RECT 3.740 3.650 4.000 3.910 ;
        RECT 6.750 3.650 7.010 3.910 ;
        RECT 3.740 0.710 4.000 0.970 ;
        RECT 6.750 0.710 7.010 0.970 ;
      LAYER met2 ;
        RECT 3.730 0.680 4.010 6.460 ;
        RECT 6.740 0.680 7.020 6.880 ;
    END
  END VSS
  PIN VDD
    ANTENNADIFFAREA 4.688600 ;
    PORT
      LAYER nwell ;
        RECT 5.160 7.560 11.180 15.120 ;
        RECT 8.600 0.000 11.180 7.560 ;
      LAYER li1 ;
        RECT 5.895 11.255 6.145 14.785 ;
        RECT 6.755 11.255 7.005 14.785 ;
        RECT 7.615 11.255 7.865 14.785 ;
        RECT 9.765 13.775 10.015 14.785 ;
        RECT 6.325 7.895 6.575 8.905 ;
        RECT 7.185 7.895 7.435 8.905 ;
        RECT 9.335 7.895 9.585 11.425 ;
        RECT 10.195 7.895 10.445 11.425 ;
        RECT 9.335 3.695 9.585 7.225 ;
        RECT 10.195 3.695 10.445 7.225 ;
        RECT 9.765 0.335 10.015 1.345 ;
      LAYER mcon ;
        RECT 5.935 13.775 6.105 13.945 ;
        RECT 6.795 13.775 6.965 13.945 ;
        RECT 7.655 13.775 7.825 13.945 ;
        RECT 9.805 14.195 9.975 14.365 ;
        RECT 6.365 8.315 6.535 8.485 ;
        RECT 7.225 8.315 7.395 8.485 ;
        RECT 9.375 8.315 9.545 8.485 ;
        RECT 10.235 8.315 10.405 8.485 ;
        RECT 9.375 6.635 9.545 6.805 ;
        RECT 10.235 6.635 10.405 6.805 ;
        RECT 9.805 0.755 9.975 0.925 ;
      LAYER met1 ;
        RECT 9.290 14.140 10.490 14.420 ;
        RECT 5.850 13.720 7.910 14.000 ;
        RECT 7.150 8.680 10.480 8.960 ;
        RECT 6.280 8.260 7.480 8.540 ;
        RECT 9.290 8.260 10.490 8.540 ;
        RECT 9.290 6.580 10.490 6.860 ;
        RECT 9.290 0.700 10.490 0.980 ;
      LAYER via ;
        RECT 10.190 14.150 10.450 14.410 ;
        RECT 7.180 13.730 7.440 13.990 ;
        RECT 7.180 8.690 7.440 8.950 ;
        RECT 10.190 8.690 10.450 8.950 ;
        RECT 7.180 8.270 7.440 8.530 ;
        RECT 10.190 8.270 10.450 8.530 ;
        RECT 10.190 6.590 10.450 6.850 ;
        RECT 10.190 0.710 10.450 0.970 ;
      LAYER met2 ;
        RECT 7.170 8.240 7.450 14.020 ;
        RECT 10.180 0.680 10.460 14.440 ;
    END
  END VDD
  PIN OUT
    ANTENNADIFFAREA 1.176000 ;
    PORT
      LAYER li1 ;
        RECT 7.185 3.695 7.435 7.225 ;
        RECT 8.045 7.055 8.295 8.065 ;
        RECT 9.765 7.895 10.015 11.425 ;
      LAYER mcon ;
        RECT 8.085 7.895 8.255 8.065 ;
        RECT 9.805 7.895 9.975 8.065 ;
        RECT 7.225 7.055 7.395 7.225 ;
        RECT 8.085 7.055 8.255 7.225 ;
      LAYER met1 ;
        RECT 8.000 7.840 10.060 8.120 ;
        RECT 7.140 7.000 8.340 7.280 ;
    END
  END OUT
  PIN INN
    ANTENNAGATEAREA 0.630000 ;
    PORT
      LAYER li1 ;
        RECT 1.165 9.995 1.415 11.005 ;
      LAYER mcon ;
        RECT 1.205 10.415 1.375 10.585 ;
      LAYER met1 ;
        RECT 0.260 10.360 1.460 10.640 ;
    END
  END INN
  PIN INP
    ANTENNAGATEAREA 0.630000 ;
    PORT
      LAYER li1 ;
        RECT 3.745 9.995 3.995 11.005 ;
      LAYER mcon ;
        RECT 3.785 10.415 3.955 10.585 ;
      LAYER met1 ;
        RECT 3.700 10.360 4.900 10.640 ;
    END
  END INP
  OBS
      LAYER pwell ;
        RECT 0.605 11.105 1.975 13.465 ;
        RECT 3.185 11.105 4.555 13.465 ;
        RECT 1.075 7.710 1.505 9.090 ;
        RECT 3.655 7.710 4.085 9.090 ;
        RECT 3.185 3.545 5.415 5.905 ;
        RECT 6.625 3.545 7.995 5.905 ;
      LAYER li1 ;
        RECT 0.735 11.255 0.985 14.785 ;
        RECT 1.165 11.255 1.415 14.785 ;
        RECT 1.595 11.255 1.845 14.785 ;
        RECT 3.315 11.255 3.565 14.785 ;
        RECT 3.745 11.255 3.995 14.785 ;
        RECT 4.175 11.255 4.425 14.785 ;
        RECT 4.605 14.615 4.855 15.205 ;
        RECT 6.325 11.255 6.575 14.785 ;
        RECT 7.185 11.255 7.435 14.785 ;
        RECT 9.765 11.675 10.015 12.685 ;
        RECT 6.325 9.995 6.575 11.005 ;
        RECT 7.185 9.995 7.435 11.005 ;
        RECT 1.165 7.895 1.415 8.905 ;
        RECT 3.745 7.895 3.995 8.905 ;
        RECT 3.745 3.695 3.995 7.225 ;
        RECT 4.605 3.695 4.855 7.225 ;
        RECT 9.765 3.695 10.015 7.225 ;
        RECT 3.745 2.435 3.995 3.445 ;
        RECT 4.605 2.435 4.855 3.445 ;
        RECT 6.325 2.855 6.575 3.445 ;
        RECT 7.185 2.435 7.435 3.445 ;
        RECT 9.765 2.435 10.015 3.445 ;
      LAYER mcon ;
        RECT 4.645 15.035 4.815 15.205 ;
        RECT 0.775 14.195 0.945 14.365 ;
        RECT 1.205 14.615 1.375 14.785 ;
        RECT 1.635 14.195 1.805 14.365 ;
        RECT 3.355 14.195 3.525 14.365 ;
        RECT 3.785 14.615 3.955 14.785 ;
        RECT 4.645 14.615 4.815 14.785 ;
        RECT 6.365 14.615 6.535 14.785 ;
        RECT 4.215 14.195 4.385 14.365 ;
        RECT 7.225 14.195 7.395 14.365 ;
        RECT 9.805 12.095 9.975 12.265 ;
        RECT 6.365 10.415 6.535 10.585 ;
        RECT 7.225 10.415 7.395 10.585 ;
        RECT 1.205 8.315 1.375 8.485 ;
        RECT 3.785 8.315 3.955 8.485 ;
        RECT 3.785 6.635 3.955 6.805 ;
        RECT 4.645 7.055 4.815 7.225 ;
        RECT 9.805 7.055 9.975 7.225 ;
        RECT 3.785 2.855 3.955 3.025 ;
        RECT 4.645 2.855 4.815 3.025 ;
        RECT 6.365 3.275 6.535 3.445 ;
        RECT 6.365 2.855 6.535 3.025 ;
        RECT 7.225 2.855 7.395 3.025 ;
        RECT 9.805 2.855 9.975 3.025 ;
      LAYER met1 ;
        RECT 4.560 14.980 6.180 15.260 ;
        RECT 0.260 14.560 3.170 14.840 ;
        RECT 3.700 14.560 4.900 14.840 ;
        RECT 5.420 14.560 6.620 14.840 ;
        RECT 0.690 14.140 1.890 14.420 ;
        RECT 3.270 14.140 4.470 14.420 ;
        RECT 5.860 14.140 7.900 14.420 ;
        RECT 7.580 12.040 10.060 12.320 ;
        RECT 6.280 10.360 7.480 10.640 ;
        RECT 1.560 9.520 3.600 9.800 ;
        RECT 0.690 8.260 1.890 8.540 ;
        RECT 3.270 8.260 4.470 8.540 ;
        RECT 4.560 7.000 5.760 7.280 ;
        RECT 8.860 7.000 10.060 7.280 ;
        RECT 3.280 6.580 4.900 6.860 ;
        RECT 4.570 3.220 6.620 3.500 ;
        RECT 8.010 3.220 10.050 3.500 ;
        RECT 3.700 2.800 4.900 3.080 ;
        RECT 6.280 2.800 8.340 3.080 ;
        RECT 8.860 2.800 10.060 3.080 ;
      LAYER via ;
        RECT 5.890 14.990 6.150 15.250 ;
        RECT 2.880 14.570 3.140 14.830 ;
        RECT 6.320 14.570 6.580 14.830 ;
        RECT 1.590 14.150 1.850 14.410 ;
        RECT 3.310 14.150 3.570 14.410 ;
        RECT 5.890 14.150 6.150 14.410 ;
        RECT 7.610 14.150 7.870 14.410 ;
        RECT 7.610 12.050 7.870 12.310 ;
        RECT 6.320 10.370 6.580 10.630 ;
        RECT 1.590 9.530 1.850 9.790 ;
        RECT 3.310 9.530 3.570 9.790 ;
        RECT 1.590 8.270 1.850 8.530 ;
        RECT 3.310 8.270 3.570 8.530 ;
        RECT 4.600 7.010 4.860 7.270 ;
        RECT 9.760 7.010 10.020 7.270 ;
        RECT 3.310 6.590 3.570 6.850 ;
        RECT 4.600 3.230 4.860 3.490 ;
        RECT 8.040 3.230 8.300 3.490 ;
        RECT 9.760 3.230 10.020 3.490 ;
        RECT 4.600 2.810 4.860 3.070 ;
        RECT 8.040 2.810 8.300 3.070 ;
        RECT 9.760 2.810 10.020 3.070 ;
      LAYER met2 ;
        RECT 1.580 8.240 1.860 14.440 ;
        RECT 2.870 13.675 3.150 14.860 ;
        RECT 3.300 6.560 3.580 14.440 ;
        RECT 5.880 14.120 6.160 15.280 ;
        RECT 6.310 10.340 6.590 14.860 ;
        RECT 7.600 12.020 7.880 14.440 ;
        RECT 4.590 2.780 4.870 7.300 ;
        RECT 8.030 2.780 8.310 3.520 ;
        RECT 9.750 2.780 10.030 7.300 ;
      LAYER via2 ;
        RECT 2.870 13.720 3.150 14.000 ;
        RECT 6.310 13.720 6.590 14.000 ;
      LAYER met3 ;
        RECT 2.845 13.460 6.615 14.260 ;
  END
END ADC_1BIT
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ADC_1BIT
  CLASS BLOCK ;
  FOREIGN ADC_1BIT ;
  ORIGIN 0.590 0.590 ;
  SIZE 13.020 BY 15.710 ;
  PIN VSS
    ANTENNADIFFAREA 3.385200 ;
    PORT
      LAYER pwell ;
        RECT 6.235 13.590 7.525 14.970 ;
        RECT 9.675 13.590 10.105 14.970 ;
      LAYER li1 ;
        RECT 6.325 13.775 6.575 14.785 ;
        RECT 7.185 13.775 7.435 14.785 ;
        RECT 9.765 13.775 10.015 14.785 ;
        RECT 5.895 7.895 6.145 11.425 ;
        RECT 6.755 7.895 7.005 11.425 ;
        RECT 7.615 7.895 7.865 11.425 ;
        RECT 9.335 7.895 9.585 11.425 ;
        RECT 10.195 7.895 10.445 11.425 ;
      LAYER mcon ;
        RECT 6.365 14.195 6.535 14.365 ;
        RECT 7.225 14.195 7.395 14.365 ;
        RECT 9.805 14.195 9.975 14.365 ;
        RECT 5.935 8.735 6.105 8.905 ;
        RECT 6.795 8.735 6.965 8.905 ;
        RECT 7.655 8.735 7.825 8.905 ;
        RECT 9.375 8.315 9.545 8.485 ;
        RECT 10.235 8.315 10.405 8.485 ;
      LAYER met1 ;
        RECT 6.280 14.140 7.480 14.420 ;
        RECT 9.290 14.140 10.490 14.420 ;
        RECT 5.850 8.680 7.910 8.960 ;
        RECT 9.290 8.260 10.490 8.540 ;
      LAYER via ;
        RECT 6.320 14.150 6.580 14.410 ;
        RECT 10.190 14.150 10.450 14.410 ;
        RECT 6.320 8.690 6.580 8.950 ;
        RECT 10.190 8.270 10.450 8.530 ;
      LAYER met2 ;
        RECT 6.310 8.635 6.590 14.440 ;
        RECT 10.180 8.240 10.460 14.440 ;
      LAYER via2 ;
        RECT 6.310 8.680 6.590 8.960 ;
        RECT 10.180 8.680 10.460 8.960 ;
      LAYER met3 ;
        RECT -0.400 8.420 12.240 9.220 ;
      LAYER via3 ;
        RECT 11.680 8.660 12.000 8.980 ;
      LAYER met4 ;
        RECT 11.250 -0.590 12.430 9.410 ;
    END
  END VSS
  PIN VDD
    ANTENNADIFFAREA 4.688600 ;
    PORT
      LAYER nwell ;
        RECT 2.580 7.560 5.160 15.120 ;
        RECT 0.000 0.000 3.440 7.560 ;
        RECT 8.600 0.000 11.180 7.560 ;
      LAYER li1 ;
        RECT 3.745 13.775 3.995 14.785 ;
        RECT 3.315 7.895 3.565 11.425 ;
        RECT 4.175 7.895 4.425 11.425 ;
        RECT 1.165 6.215 1.415 7.225 ;
        RECT 2.025 6.215 2.275 7.225 ;
        RECT 0.735 0.335 0.985 3.865 ;
        RECT 1.595 0.335 1.845 3.865 ;
        RECT 2.455 0.335 2.705 3.865 ;
        RECT 9.335 3.695 9.585 7.225 ;
        RECT 10.195 3.695 10.445 7.225 ;
        RECT 9.765 0.335 10.015 1.345 ;
      LAYER mcon ;
        RECT 3.785 14.195 3.955 14.365 ;
        RECT 3.355 8.315 3.525 8.485 ;
        RECT 4.215 8.315 4.385 8.485 ;
        RECT 1.205 6.635 1.375 6.805 ;
        RECT 2.065 6.635 2.235 6.805 ;
        RECT 9.375 6.635 9.545 6.805 ;
        RECT 0.775 1.175 0.945 1.345 ;
        RECT 1.635 1.175 1.805 1.345 ;
        RECT 10.235 6.635 10.405 6.805 ;
        RECT 2.495 1.175 2.665 1.345 ;
        RECT 9.805 0.755 9.975 0.925 ;
      LAYER met1 ;
        RECT 3.270 14.140 4.470 14.420 ;
        RECT 4.140 8.680 4.890 8.960 ;
        RECT 3.270 8.260 4.470 8.540 ;
        RECT 1.120 6.580 2.320 6.860 ;
        RECT 9.290 6.580 10.490 6.860 ;
        RECT 0.690 1.120 2.750 1.400 ;
        RECT 9.290 0.700 10.490 0.980 ;
        RECT 9.730 0.280 10.480 0.560 ;
      LAYER via ;
        RECT 4.170 14.150 4.430 14.410 ;
        RECT 4.170 8.690 4.430 8.950 ;
        RECT 4.600 8.690 4.860 8.950 ;
        RECT 4.170 8.270 4.430 8.530 ;
        RECT 1.160 6.590 1.420 6.850 ;
        RECT 10.190 6.590 10.450 6.850 ;
        RECT 1.160 1.130 1.420 1.390 ;
        RECT 10.190 0.710 10.450 0.970 ;
        RECT 9.760 0.290 10.020 0.550 ;
        RECT 10.190 0.290 10.450 0.550 ;
      LAYER met2 ;
        RECT 4.160 8.240 4.440 14.440 ;
        RECT 1.150 -0.185 1.430 6.880 ;
        RECT 4.590 -0.185 4.870 8.980 ;
        RECT 9.750 -0.185 10.030 0.580 ;
        RECT 10.180 0.260 10.460 6.880 ;
      LAYER via2 ;
        RECT 1.150 -0.140 1.430 0.140 ;
        RECT 4.590 -0.140 4.870 0.140 ;
        RECT 9.750 -0.140 10.030 0.140 ;
      LAYER met3 ;
        RECT -0.400 -0.400 12.240 0.400 ;
      LAYER via3 ;
        RECT -0.160 -0.160 0.160 0.160 ;
      LAYER met4 ;
        RECT -0.590 -0.590 0.590 9.410 ;
    END
  END VDD
  PIN OUT
    ANTENNADIFFAREA 1.176000 ;
    PORT
      LAYER li1 ;
        RECT 9.765 7.895 10.015 11.425 ;
        RECT 9.765 3.695 10.015 7.225 ;
      LAYER mcon ;
        RECT 9.805 7.895 9.975 8.065 ;
        RECT 9.805 7.055 9.975 7.225 ;
      LAYER met1 ;
        RECT 8.860 7.840 10.060 8.120 ;
        RECT 8.860 7.000 10.060 7.280 ;
      LAYER via ;
        RECT 9.330 7.850 9.590 8.110 ;
        RECT 9.330 7.010 9.590 7.270 ;
      LAYER met2 ;
        RECT 9.320 6.980 9.600 8.140 ;
    END
  END OUT
  PIN INN
    ANTENNAGATEAREA 0.630000 ;
    PORT
      LAYER li1 ;
        RECT 4.605 4.115 4.855 5.125 ;
      LAYER mcon ;
        RECT 4.645 4.535 4.815 4.705 ;
      LAYER met1 ;
        RECT 3.700 4.480 4.900 4.760 ;
    END
  END INN
  PIN INP
    ANTENNAGATEAREA 0.630000 ;
    PORT
      LAYER li1 ;
        RECT 7.185 4.115 7.435 5.125 ;
      LAYER mcon ;
        RECT 7.225 4.535 7.395 4.705 ;
      LAYER met1 ;
        RECT 7.140 4.480 8.340 4.760 ;
    END
  END INP
  OBS
      LAYER pwell ;
        RECT 5.765 9.215 7.995 11.575 ;
        RECT 9.205 9.215 10.575 11.575 ;
        RECT 4.515 6.030 4.945 7.410 ;
        RECT 7.095 6.030 7.525 7.410 ;
        RECT 4.045 1.655 5.415 4.015 ;
        RECT 6.625 1.655 7.995 4.015 ;
      LAYER li1 ;
        RECT 3.745 11.675 3.995 12.685 ;
        RECT 6.325 11.675 6.575 12.685 ;
        RECT 7.185 11.675 7.435 12.685 ;
        RECT 8.475 11.675 8.725 12.265 ;
        RECT 9.765 11.675 10.015 12.685 ;
        RECT 3.745 7.895 3.995 11.425 ;
        RECT 6.325 7.895 6.575 11.425 ;
        RECT 7.185 7.895 7.435 11.425 ;
        RECT 4.605 6.215 4.855 7.225 ;
        RECT 7.185 6.215 7.435 7.225 ;
        RECT 1.165 4.115 1.415 5.125 ;
        RECT 2.025 4.115 2.275 5.125 ;
        RECT 1.165 0.335 1.415 3.865 ;
        RECT 2.025 0.335 2.275 3.865 ;
        RECT 3.315 0.755 3.565 1.345 ;
        RECT 4.175 0.335 4.425 3.865 ;
        RECT 4.605 0.335 4.855 3.865 ;
        RECT 5.035 0.335 5.285 3.865 ;
        RECT 6.325 0.335 6.575 1.345 ;
        RECT 6.755 0.335 7.005 3.865 ;
        RECT 7.185 0.335 7.435 3.865 ;
        RECT 7.615 0.335 7.865 3.865 ;
        RECT 8.045 0.335 8.295 3.025 ;
        RECT 9.765 2.435 10.015 3.445 ;
      LAYER mcon ;
        RECT 3.785 12.095 3.955 12.265 ;
        RECT 6.365 12.095 6.535 12.265 ;
        RECT 7.225 12.095 7.395 12.265 ;
        RECT 8.515 12.095 8.685 12.265 ;
        RECT 8.515 11.675 8.685 11.845 ;
        RECT 9.805 12.095 9.975 12.265 ;
        RECT 3.785 7.895 3.955 8.065 ;
        RECT 6.365 8.315 6.535 8.485 ;
        RECT 7.225 7.895 7.395 8.065 ;
        RECT 4.645 6.635 4.815 6.805 ;
        RECT 7.225 6.635 7.395 6.805 ;
        RECT 1.205 4.535 1.375 4.705 ;
        RECT 2.065 4.535 2.235 4.705 ;
        RECT 1.205 0.755 1.375 0.925 ;
        RECT 3.355 1.175 3.525 1.345 ;
        RECT 3.355 0.755 3.525 0.925 ;
        RECT 4.215 0.755 4.385 0.925 ;
        RECT 2.065 0.335 2.235 0.505 ;
        RECT 4.645 0.335 4.815 0.505 ;
        RECT 5.075 0.755 5.245 0.925 ;
        RECT 6.365 1.175 6.535 1.345 ;
        RECT 6.365 0.335 6.535 0.505 ;
        RECT 6.795 0.755 6.965 0.925 ;
        RECT 7.225 0.335 7.395 0.505 ;
        RECT 7.655 0.755 7.825 0.925 ;
        RECT 8.085 2.855 8.255 3.025 ;
        RECT 9.805 2.855 9.975 3.025 ;
        RECT 8.085 0.335 8.255 0.505 ;
      LAYER met1 ;
        RECT 2.840 12.040 4.040 12.320 ;
        RECT 6.280 12.040 7.480 12.320 ;
        RECT 8.430 12.040 10.060 12.320 ;
        RECT 3.710 11.620 8.770 11.900 ;
        RECT 6.280 8.260 7.480 8.540 ;
        RECT 2.840 7.840 4.040 8.120 ;
        RECT 7.140 7.840 8.340 8.120 ;
        RECT 4.130 6.580 5.330 6.860 ;
        RECT 6.710 6.580 7.910 6.860 ;
        RECT 5.000 5.320 7.040 5.600 ;
        RECT 1.120 4.480 2.320 4.760 ;
        RECT 8.000 2.800 10.060 3.080 ;
        RECT 3.270 1.120 6.620 1.400 ;
        RECT 1.120 0.700 3.610 0.980 ;
        RECT 4.130 0.700 5.330 0.980 ;
        RECT 6.710 0.700 7.910 0.980 ;
        RECT 1.980 0.280 3.180 0.560 ;
        RECT 3.700 0.280 4.900 0.560 ;
        RECT 6.280 0.280 8.340 0.560 ;
      LAYER via ;
        RECT 3.740 12.050 4.000 12.310 ;
        RECT 7.180 12.050 7.440 12.310 ;
        RECT 3.740 11.630 4.000 11.890 ;
        RECT 7.180 11.630 7.440 11.890 ;
        RECT 6.750 8.270 7.010 8.530 ;
        RECT 3.740 7.850 4.000 8.110 ;
        RECT 7.180 7.850 7.440 8.110 ;
        RECT 5.030 6.590 5.290 6.850 ;
        RECT 6.750 6.590 7.010 6.850 ;
        RECT 5.030 5.330 5.290 5.590 ;
        RECT 6.750 5.330 7.010 5.590 ;
        RECT 2.020 4.490 2.280 4.750 ;
        RECT 5.030 0.710 5.290 0.970 ;
        RECT 6.750 0.710 7.010 0.970 ;
        RECT 2.020 0.290 2.280 0.550 ;
        RECT 3.740 0.290 4.000 0.550 ;
      LAYER met2 ;
        RECT 3.730 7.820 4.010 12.340 ;
        RECT 2.010 0.260 2.290 4.780 ;
        RECT 3.730 0.260 4.010 1.445 ;
        RECT 5.020 0.680 5.300 6.880 ;
        RECT 6.740 0.680 7.020 8.560 ;
        RECT 7.170 7.820 7.450 12.340 ;
      LAYER via2 ;
        RECT 2.010 1.120 2.290 1.400 ;
        RECT 3.730 1.120 4.010 1.400 ;
      LAYER met3 ;
        RECT 1.985 0.860 4.035 1.660 ;
  END
END ADC_1BIT
END LIBRARY


magic
tech sky130A
timestamp 1676315893
<< end >>

module msvsd4bituc (INN,
    OUT,
    \r_VSS(0) ,
    \r_VSS(1) ,
    \r_VSS(2) ,
    \r_VDD(0) ,
    \r_VDD(1) ,
    \r_VDD(2) );
 input INN;
 output OUT;
 input \r_VSS(0) ;
 input \r_VSS(1) ;
 input \r_VSS(2) ;
 input \r_VDD(0) ;
 input \r_VDD(1) ;
 input \r_VDD(2) ;

 wire ring_adc;
 wire r_VSS;
 wire r_VDD;

 ADC_1BIT ADC_1BIT (.OUT(OUT),
    .INN(INN),
    .INP(ring_adc));
 RING_OSCILLATOR RING_OSCILLATOR (.INP(ring_adc));
 sky130_fd_sc_hd__decap_4 PHY_0 ();
 sky130_fd_sc_hd__decap_4 PHY_1 ();
 sky130_fd_sc_hd__decap_4 PHY_2 ();
 sky130_fd_sc_hd__decap_4 PHY_3 ();
 sky130_fd_sc_hd__decap_4 PHY_4 ();
 sky130_fd_sc_hd__decap_4 PHY_5 ();
 sky130_fd_sc_hd__decap_4 PHY_6 ();
 sky130_fd_sc_hd__decap_4 PHY_7 ();
 sky130_fd_sc_hd__decap_4 PHY_8 ();
 sky130_fd_sc_hd__decap_4 PHY_9 ();
 sky130_fd_sc_hd__decap_4 PHY_10 ();
 sky130_fd_sc_hd__decap_4 PHY_11 ();
 sky130_fd_sc_hd__decap_4 PHY_12 ();
 sky130_fd_sc_hd__decap_4 PHY_13 ();
 sky130_fd_sc_hd__decap_4 PHY_14 ();
 sky130_fd_sc_hd__decap_4 PHY_15 ();
 sky130_fd_sc_hd__decap_4 PHY_16 ();
 sky130_fd_sc_hd__decap_4 PHY_17 ();
 sky130_fd_sc_hd__decap_4 PHY_18 ();
 sky130_fd_sc_hd__decap_4 PHY_19 ();
 sky130_fd_sc_hd__decap_4 PHY_20 ();
 sky130_fd_sc_hd__decap_4 PHY_21 ();
 sky130_fd_sc_hd__decap_4 PHY_22 ();
 sky130_fd_sc_hd__decap_4 PHY_23 ();
 sky130_fd_sc_hd__decap_4 PHY_24 ();
 sky130_fd_sc_hd__decap_4 PHY_25 ();
 sky130_fd_sc_hd__decap_4 PHY_26 ();
 sky130_fd_sc_hd__decap_4 PHY_27 ();
 sky130_fd_sc_hd__decap_4 PHY_28 ();
 sky130_fd_sc_hd__decap_4 PHY_29 ();
 sky130_fd_sc_hd__decap_4 PHY_30 ();
 sky130_fd_sc_hd__decap_4 PHY_31 ();
 sky130_fd_sc_hd__decap_4 PHY_32 ();
 sky130_fd_sc_hd__decap_4 PHY_33 ();
 sky130_fd_sc_hd__decap_4 PHY_34 ();
 sky130_fd_sc_hd__decap_4 PHY_35 ();
 sky130_fd_sc_hd__decap_4 PHY_36 ();
 sky130_fd_sc_hd__decap_4 PHY_37 ();
 sky130_fd_sc_hd__decap_4 PHY_38 ();
 sky130_fd_sc_hd__decap_4 PHY_39 ();
 sky130_fd_sc_hd__decap_4 PHY_40 ();
 sky130_fd_sc_hd__decap_4 PHY_41 ();
 sky130_fd_sc_hd__decap_4 PHY_42 ();
 sky130_fd_sc_hd__decap_4 PHY_43 ();
 sky130_fd_sc_hd__decap_4 PHY_44 ();
 sky130_fd_sc_hd__decap_4 PHY_45 ();
 sky130_fd_sc_hd__decap_4 PHY_46 ();
 sky130_fd_sc_hd__decap_4 PHY_47 ();
 sky130_fd_sc_hd__decap_4 PHY_48 ();
 sky130_fd_sc_hd__decap_4 PHY_49 ();
 sky130_fd_sc_hd__decap_4 PHY_50 ();
 sky130_fd_sc_hd__decap_4 PHY_51 ();
 sky130_fd_sc_hd__decap_4 PHY_52 ();
 sky130_fd_sc_hd__decap_4 PHY_53 ();
 sky130_fd_sc_hd__decap_4 PHY_54 ();
 sky130_fd_sc_hd__decap_4 PHY_55 ();
 sky130_fd_sc_hd__decap_4 PHY_56 ();
 sky130_fd_sc_hd__decap_4 PHY_57 ();
 sky130_fd_sc_hd__decap_4 PHY_58 ();
 sky130_fd_sc_hd__decap_4 PHY_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_73 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_4 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_57 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_65 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_144 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_156 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_157 ();
endmodule

module RING_OSCILLATOR(
	output INP
);

endmodule

* SPICE3 file created from FUNCTION_0.ext - technology: sky130A

** sch_path: /home/syedimaduddin/Desktop/VSD PD Research Program/Week-2/xschem/function.sch
**.subckt function
XM1 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net3 C net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net3 D net2 net2 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 Y E net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Y F net3 net3 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 Y A net4 net4 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 Y C net4 net4 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 Y E net5 net5 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 net4 B GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 net4 D GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 net5 F GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
VA A GND pulse(0 1.8 0ns 1ns 1ns 4ns 10ns)
.save i(va)
VB B GND pulse(0 1.8 0.1ns 1ns 1ns 4ns 10ns)
.save i(vb)
VC C GND pulse(0 1.8 0.2ns 1ns 1ns 4ns 10ns)
.save i(vc)
VD D GND pulse(0 1.8 0.3ns 1ns 1ns 4ns 10ns)
.save i(vd)
VE E GND pulse(0 1.8 0.4ns 1ns 1ns 4ns 10ns)
.save i(ve)
VF F GND pulse(0 1.8 0.5ns 1ns 1ns 4ns 10ns)
.save i(vf)
Vdd VDD GND 1.8
.save i(vdd)
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt



.tran 0.01n 60n
.save all


**** end user architecture code
**.ends

.GLOBAL VDD
.GLOBAL GND


.subckt NMOS_S_79666698_X5_Y1_1676686594 a_230_462# a_200_252# a_147_462#
X0 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=1.47e+12p pd=1.33e+07u as=1.7325e+12p ps=1.59e+07u w=1.05e+06u l=150000u
X1 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X2 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X3 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X4 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X5 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X6 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X7 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X8 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X9 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
C0 a_200_252# a_230_462# 0.56fF
C1 a_230_462# a_147_462# 3.74fF
C2 a_200_252# a_147_462# 3.07fF
.ends

.subckt PMOS_S_49267959_X5_Y1_1676686590_1676686592 a_230_357# a_200_252# w_0_0# VSUBS
X0 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.94e+12p pd=2.38e+07u as=3.465e+12p ps=2.85e+07u w=2.1e+06u l=150000u
X1 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X2 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X3 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X4 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X5 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X6 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X7 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X8 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X9 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
C0 w_0_0# a_200_252# 2.20fF
C1 a_230_357# a_200_252# 0.44fF
C2 a_230_357# w_0_0# 3.98fF
C3 a_230_357# VSUBS -0.16fF
C4 a_200_252# VSUBS 0.16fF
C5 w_0_0# VSUBS 5.49fF
.ends

.subckt NMOS_S_79666698_X5_Y1_1676686589_1676686592 a_230_462# a_200_252# a_147_462#
X0 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=1.47e+12p pd=1.33e+07u as=1.7325e+12p ps=1.59e+07u w=1.05e+06u l=150000u
X1 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X2 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X3 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X4 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X5 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X6 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X7 a_230_462# a_200_252# a_147_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X8 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X9 a_147_462# a_200_252# a_230_462# a_147_462# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
C0 a_200_252# a_230_462# 0.56fF
C1 a_230_462# a_147_462# 3.74fF
C2 a_200_252# a_147_462# 3.07fF
.ends

.subckt INV_61857474_0_0_1676686592 m1_570_1400# PMOS_S_49267959_X5_Y1_1676686590_1676686592_0/w_0_0#
+ m1_656_560# VSUBS
XPMOS_S_49267959_X5_Y1_1676686590_1676686592_0 m1_570_1400# m1_656_560# PMOS_S_49267959_X5_Y1_1676686590_1676686592_0/w_0_0#
+ VSUBS PMOS_S_49267959_X5_Y1_1676686590_1676686592
XNMOS_S_79666698_X5_Y1_1676686589_1676686592_0 m1_570_1400# m1_656_560# VSUBS NMOS_S_79666698_X5_Y1_1676686589_1676686592
C0 m1_570_1400# m1_656_560# 0.31fF
C1 PMOS_S_49267959_X5_Y1_1676686590_1676686592_0/w_0_0# m1_656_560# 0.41fF
C2 PMOS_S_49267959_X5_Y1_1676686590_1676686592_0/w_0_0# m1_570_1400# 0.05fF
C3 m1_570_1400# VSUBS 3.26fF
C4 m1_656_560# VSUBS 3.70fF
C5 PMOS_S_49267959_X5_Y1_1676686590_1676686592_0/w_0_0# VSUBS 5.63fF
.ends

.subckt DP_PMOS_34936022_X5_Y1_1676686593 a_372_252# a_230_357# a_200_252# a_402_357#
+ w_0_0# VSUBS
X0 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.94e+12p pd=2.38e+07u as=6.405e+12p ps=5.23e+07u w=2.1e+06u l=150000u
X1 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X2 a_402_357# a_372_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.94e+12p pd=2.38e+07u as=0p ps=0u w=2.1e+06u l=150000u
X3 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X4 a_402_357# a_372_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X5 a_402_357# a_372_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X6 w_0_0# a_372_252# a_402_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X7 w_0_0# a_372_252# a_402_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X8 a_402_357# a_372_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X9 a_402_357# a_372_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X10 w_0_0# a_372_252# a_402_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X11 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X12 w_0_0# a_372_252# a_402_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X13 w_0_0# a_372_252# a_402_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X14 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X15 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X16 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X17 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X18 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X19 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
C0 a_230_357# a_200_252# 0.45fF
C1 a_372_252# w_0_0# 2.29fF
C2 a_200_252# w_0_0# 2.35fF
C3 a_372_252# a_402_357# 0.43fF
C4 a_200_252# a_402_357# 0.05fF
C5 a_372_252# a_200_252# 2.09fF
C6 a_230_357# w_0_0# 3.48fF
C7 a_230_357# a_402_357# 0.88fF
C8 a_372_252# a_230_357# 0.02fF
C9 w_0_0# a_402_357# 4.75fF
C10 a_402_357# VSUBS -0.30fF
C11 a_230_357# VSUBS -0.24fF
C12 a_372_252# VSUBS 0.06fF
C13 a_200_252# VSUBS -0.14fF
C14 w_0_0# VSUBS 8.10fF
.ends

.subckt PMOS_S_49267959_X5_Y1_1676686595 a_230_357# a_200_252# w_0_0# VSUBS
X0 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.94e+12p pd=2.38e+07u as=3.465e+12p ps=2.85e+07u w=2.1e+06u l=150000u
X1 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X2 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X3 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X4 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X5 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X6 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X7 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X8 a_230_357# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
X9 w_0_0# a_200_252# a_230_357# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.1e+06u l=150000u
C0 a_230_357# w_0_0# 3.98fF
C1 a_200_252# w_0_0# 2.20fF
C2 a_230_357# a_200_252# 0.44fF
C3 a_230_357# VSUBS -0.16fF
C4 a_200_252# VSUBS 0.16fF
C5 w_0_0# VSUBS 5.49fF
.ends

.subckt FUNCTION_0 Y A B C D E F VDD GND
XNMOS_S_79666698_X5_Y1_1676686594_0 Y C GND NMOS_S_79666698_X5_Y1_1676686594
XNMOS_S_79666698_X5_Y1_1676686594_1 Y A GND NMOS_S_79666698_X5_Y1_1676686594
XNMOS_S_79666698_X5_Y1_1676686594_2 GND m1_946_2408# GND NMOS_S_79666698_X5_Y1_1676686594
XNMOS_S_79666698_X5_Y1_1676686594_3 GND D GND NMOS_S_79666698_X5_Y1_1676686594
XNMOS_S_79666698_X5_Y1_1676686594_4 GND m1_2720_560# GND NMOS_S_79666698_X5_Y1_1676686594
XINV_61857474_0_0_1676686592_0 Y w_3328_1530# E GND INV_61857474_0_0_1676686592
XDP_PMOS_34936022_X5_Y1_1676686593_0 m1_2720_560# w_3328_1530# A w_3328_1530# VDD
+ GND DP_PMOS_34936022_X5_Y1_1676686593
XPMOS_S_49267959_X5_Y1_1676686595_0 Y m1_946_2408# w_3328_1530# GND PMOS_S_49267959_X5_Y1_1676686595
XPMOS_S_49267959_X5_Y1_1676686595_1 w_3328_1530# D w_3328_1530# GND PMOS_S_49267959_X5_Y1_1676686595
XPMOS_S_49267959_X5_Y1_1676686595_2 w_3328_1530# C w_3328_1530# GND PMOS_S_49267959_X5_Y1_1676686595
C0 m1_946_2408# C 0.29fF
C1 A C 0.33fF
C2 VDD C 0.02fF
C3 E m1_946_2408# 0.01fF
C4 A m1_946_2408# 0.15fF
C5 VDD m1_946_2408# 0.03fF
C6 D Y 0.06fF
C7 VDD A 0.35fF
C8 D w_3328_1530# 1.11fF
C9 D B 0.04fF
C10 Y w_3328_1530# 3.02fF
C11 B Y 0.05fF
C12 B w_3328_1530# 0.76fF
C13 D m1_2720_560# 0.18fF
C14 m1_2720_560# Y 0.12fF
C15 m1_2720_560# w_3328_1530# 0.90fF
C16 D C 0.07fF
C17 Y C 0.16fF
C18 w_3328_1530# C 1.33fF
C19 B C 0.01fF
C20 D E 0.03fF
C21 Y E 0.02fF
C22 D m1_946_2408# 0.27fF
C23 m1_2720_560# C 0.01fF
C24 E w_3328_1530# 0.08fF
C25 Y m1_946_2408# 0.34fF
C26 B E 0.03fF
C27 D A 0.01fF
C28 D VDD 0.02fF
C29 Y A 0.34fF
C30 m1_946_2408# w_3328_1530# 0.83fF
C31 B m1_946_2408# 0.00fF
C32 A w_3328_1530# 1.49fF
C33 VDD w_3328_1530# 0.16fF
C34 B A 0.04fF
C35 m1_2720_560# m1_946_2408# 0.15fF
C36 m1_2720_560# A 0.33fF
C37 VDD m1_2720_560# 0.35fF
C38 B GND 0.32fF **FLOATING
C39 Y GND 9.54fF
C40 w_3328_1530# GND 21.22fF
C41 A GND 2.79fF
C42 C GND 2.94fF
C43 D GND 3.46fF
C44 m1_946_2408# GND 4.40fF
C45 VDD GND 8.48fF
C46 E GND 3.22fF
C47 m1_2720_560# GND 3.97fF
.ends

